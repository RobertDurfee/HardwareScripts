#INCLUDES

module Synth(
  input bit clk,
  #INPUTS,
  output #OUTPUT_TYPE out
);

  assign out = #FUNCTION_CALL;

endmodule
