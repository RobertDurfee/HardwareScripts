module $CELL_NAME(
  $INPUTS,
  $OUTPUTS
);

  $OUTPUT_FUNCTIONS;

endmodule
